-----------------------------------------------------------------------
--
--  test bench para o gerado de padr�es
--
--  Fernando Moraes
-----------------------------------------------------------------------
library ieee;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_1164.all;


entity user_logic_tb is
end user_logic_tb;

architecture TB_ARCHITECTURE of user_logic_tb is         


begin
  
         
end TB_ARCHITECTURE;
